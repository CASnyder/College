--***************************************************************
--VHDL CODE FOR SECTION 4.2(A)
-- Authors: C. A. Snyder
--				B. Rutledge
--				M. Bbela 	
--			
-- File: enhanced_prio.vhd
--
-- Design units:
--
-- ENTITY enhanced_prio
-- ARCHITECTURE prio_arch
-- Purpose:  
-- Inputs: r: 10 bit input request
-- Outputs: fst: 4 bit, binary code of the highest priority request
--				snd: 4 bit, binary code of the second-highest priority request 
-- 
-- Library/Package:
-- ieee.std_logic_1164: to use std_logic
--
-- Software/Version:
-- Simulated by: Altera Quartus v13.0.1
-- Synthesized by: Altera Quartus v13.0.1
--
-- Revision History
-- Version 1.0:
-- Date: 9/21/2015
-- Comments: Original
--
--*************************************************************** 
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;	
ENTITY enhanced_prio IS 
	PORT(
		r: IN std_logic_vector(9 DOWNTO 0);
		fst, snd: OUT std_logic_vector(3 DOWNTO 0)
	);
END enhanced_prio;
ARCHITECTURE table_arch OF enhanced_prio IS
		SIGNAL both: std_logic_vector(7 downto 0);
BEGIN
	WITH r SELECT
		both <= 
"11111111" when "0000000000",
"00001111" when "0000000001",
"00011111" when "0000000010",
"00010000" when "0000000011",
"00101111" when "0000000100",
"00100000" when "0000000101",
"00100001" when "0000000110",
"00100001" when "0000000111",
"00111111" when "0000001000",
"00110000" when "0000001001",
"00110001" when "0000001010",
"00110001" when "0000001011",
"00110010" when "0000001100",
"00110010" when "0000001101",
"00110010" when "0000001110",
"00110010" when "0000001111",
"01001111" when "0000010000",
"01000000" when "0000010001",
"01000001" when "0000010010",
"01000001" when "0000010011",
"01000010" when "0000010100",
"01000010" when "0000010101",
"01000010" when "0000010110",
"01000010" when "0000010111",
"01000011" when "0000011000",
"01000011" when "0000011001",
"01000011" when "0000011010",
"01000011" when "0000011011",
"01000011" when "0000011100",
"01000011" when "0000011101",
"01000011" when "0000011110",
"01000011" when "0000011111",
"01011111" when "0000100000",
"01010000" when "0000100001",
"01010001" when "0000100010",
"01010001" when "0000100011",
"01010010" when "0000100100",
"01010010" when "0000100101",
"01010010" when "0000100110",
"01010010" when "0000100111",
"01010011" when "0000101000",
"01010011" when "0000101001",
"01010011" when "0000101010",
"01010011" when "0000101011",
"01010011" when "0000101100",
"01010011" when "0000101101",
"01010011" when "0000101110",
"01010011" when "0000101111",
"01010100" when "0000110000",
"01010100" when "0000110001",
"01010100" when "0000110010",
"01010100" when "0000110011",
"01010100" when "0000110100",
"01010100" when "0000110101",
"01010100" when "0000110110",
"01010100" when "0000110111",
"01010100" when "0000111000",
"01010100" when "0000111001",
"01010100" when "0000111010",
"01010100" when "0000111011",
"01010100" when "0000111100",
"01010100" when "0000111101",
"01010100" when "0000111110",
"01010100" when "0000111111",
"01101111" when "0001000000",
"01100000" when "0001000001",
"01100001" when "0001000010",
"01100001" when "0001000011",
"01100010" when "0001000100",
"01100010" when "0001000101",
"01100010" when "0001000110",
"01100010" when "0001000111",
"01100011" when "0001001000",
"01100011" when "0001001001",
"01100011" when "0001001010",
"01100011" when "0001001011",
"01100011" when "0001001100",
"01100011" when "0001001101",
"01100011" when "0001001110",
"01100011" when "0001001111",
"01100100" when "0001010000",
"01100100" when "0001010001",
"01100100" when "0001010010",
"01100100" when "0001010011",
"01100100" when "0001010100",
"01100100" when "0001010101",
"01100100" when "0001010110",
"01100100" when "0001010111",
"01100100" when "0001011000",
"01100100" when "0001011001",
"01100100" when "0001011010",
"01100100" when "0001011011",
"01100100" when "0001011100",
"01100100" when "0001011101",
"01100100" when "0001011110",
"01100100" when "0001011111",
"01100101" when "0001100000",
"01100101" when "0001100001",
"01100101" when "0001100010",
"01100101" when "0001100011",
"01100101" when "0001100100",
"01100101" when "0001100101",
"01100101" when "0001100110",
"01100101" when "0001100111",
"01100101" when "0001101000",
"01100101" when "0001101001",
"01100101" when "0001101010",
"01100101" when "0001101011",
"01100101" when "0001101100",
"01100101" when "0001101101",
"01100101" when "0001101110",
"01100101" when "0001101111",
"01100101" when "0001110000",
"01100101" when "0001110001",
"01100101" when "0001110010",
"01100101" when "0001110011",
"01100101" when "0001110100",
"01100101" when "0001110101",
"01100101" when "0001110110",
"01100101" when "0001110111",
"01100101" when "0001111000",
"01100101" when "0001111001",
"01100101" when "0001111010",
"01100101" when "0001111011",
"01100101" when "0001111100",
"01100101" when "0001111101",
"01100101" when "0001111110",
"01100101" when "0001111111",
"01111111" when "0010000000",
"01110000" when "0010000001",
"01110001" when "0010000010",
"01110001" when "0010000011",
"01110010" when "0010000100",
"01110010" when "0010000101",
"01110010" when "0010000110",
"01110010" when "0010000111",
"01110011" when "0010001000",
"01110011" when "0010001001",
"01110011" when "0010001010",
"01110011" when "0010001011",
"01110011" when "0010001100",
"01110011" when "0010001101",
"01110011" when "0010001110",
"01110011" when "0010001111",
"01110100" when "0010010000",
"01110100" when "0010010001",
"01110100" when "0010010010",
"01110100" when "0010010011",
"01110100" when "0010010100",
"01110100" when "0010010101",
"01110100" when "0010010110",
"01110100" when "0010010111",
"01110100" when "0010011000",
"01110100" when "0010011001",
"01110100" when "0010011010",
"01110100" when "0010011011",
"01110100" when "0010011100",
"01110100" when "0010011101",
"01110100" when "0010011110",
"01110100" when "0010011111",
"01110101" when "0010100000",
"01110101" when "0010100001",
"01110101" when "0010100010",
"01110101" when "0010100011",
"01110101" when "0010100100",
"01110101" when "0010100101",
"01110101" when "0010100110",
"01110101" when "0010100111",
"01110101" when "0010101000",
"01110101" when "0010101001",
"01110101" when "0010101010",
"01110101" when "0010101011",
"01110101" when "0010101100",
"01110101" when "0010101101",
"01110101" when "0010101110",
"01110101" when "0010101111",
"01110101" when "0010110000",
"01110101" when "0010110001",
"01110101" when "0010110010",
"01110101" when "0010110011",
"01110101" when "0010110100",
"01110101" when "0010110101",
"01110101" when "0010110110",
"01110101" when "0010110111",
"01110101" when "0010111000",
"01110101" when "0010111001",
"01110101" when "0010111010",
"01110101" when "0010111011",
"01110101" when "0010111100",
"01110101" when "0010111101",
"01110101" when "0010111110",
"01110101" when "0010111111",
"01110110" when "0011000000",
"01110110" when "0011000001",
"01110110" when "0011000010",
"01110110" when "0011000011",
"01110110" when "0011000100",
"01110110" when "0011000101",
"01110110" when "0011000110",
"01110110" when "0011000111",
"01110110" when "0011001000",
"01110110" when "0011001001",
"01110110" when "0011001010",
"01110110" when "0011001011",
"01110110" when "0011001100",
"01110110" when "0011001101",
"01110110" when "0011001110",
"01110110" when "0011001111",
"01110110" when "0011010000",
"01110110" when "0011010001",
"01110110" when "0011010010",
"01110110" when "0011010011",
"01110110" when "0011010100",
"01110110" when "0011010101",
"01110110" when "0011010110",
"01110110" when "0011010111",
"01110110" when "0011011000",
"01110110" when "0011011001",
"01110110" when "0011011010",
"01110110" when "0011011011",
"01110110" when "0011011100",
"01110110" when "0011011101",
"01110110" when "0011011110",
"01110110" when "0011011111",
"01110110" when "0011100000",
"01110110" when "0011100001",
"01110110" when "0011100010",
"01110110" when "0011100011",
"01110110" when "0011100100",
"01110110" when "0011100101",
"01110110" when "0011100110",
"01110110" when "0011100111",
"01110110" when "0011101000",
"01110110" when "0011101001",
"01110110" when "0011101010",
"01110110" when "0011101011",
"01110110" when "0011101100",
"01110110" when "0011101101",
"01110110" when "0011101110",
"01110110" when "0011101111",
"01110110" when "0011110000",
"01110110" when "0011110001",
"01110110" when "0011110010",
"01110110" when "0011110011",
"01110110" when "0011110100",
"01110110" when "0011110101",
"01110110" when "0011110110",
"01110110" when "0011110111",
"01110110" when "0011111000",
"01110110" when "0011111001",
"01110110" when "0011111010",
"01110110" when "0011111011",
"01110110" when "0011111100",
"01110110" when "0011111101",
"01110110" when "0011111110",
"01110110" when "0011111111",
"10001111" when "0100000000",
"10000000" when "0100000001",
"10000001" when "0100000010",
"10000001" when "0100000011",
"10000010" when "0100000100",
"10000010" when "0100000101",
"10000010" when "0100000110",
"10000010" when "0100000111",
"10000011" when "0100001000",
"10000011" when "0100001001",
"10000011" when "0100001010",
"10000011" when "0100001011",
"10000011" when "0100001100",
"10000011" when "0100001101",
"10000011" when "0100001110",
"10000011" when "0100001111",
"10000100" when "0100010000",
"10000100" when "0100010001",
"10000100" when "0100010010",
"10000100" when "0100010011",
"10000100" when "0100010100",
"10000100" when "0100010101",
"10000100" when "0100010110",
"10000100" when "0100010111",
"10000100" when "0100011000",
"10000100" when "0100011001",
"10000100" when "0100011010",
"10000100" when "0100011011",
"10000100" when "0100011100",
"10000100" when "0100011101",
"10000100" when "0100011110",
"10000100" when "0100011111",
"10000101" when "0100100000",
"10000101" when "0100100001",
"10000101" when "0100100010",
"10000101" when "0100100011",
"10000101" when "0100100100",
"10000101" when "0100100101",
"10000101" when "0100100110",
"10000101" when "0100100111",
"10000101" when "0100101000",
"10000101" when "0100101001",
"10000101" when "0100101010",
"10000101" when "0100101011",
"10000101" when "0100101100",
"10000101" when "0100101101",
"10000101" when "0100101110",
"10000101" when "0100101111",
"10000101" when "0100110000",
"10000101" when "0100110001",
"10000101" when "0100110010",
"10000101" when "0100110011",
"10000101" when "0100110100",
"10000101" when "0100110101",
"10000101" when "0100110110",
"10000101" when "0100110111",
"10000101" when "0100111000",
"10000101" when "0100111001",
"10000101" when "0100111010",
"10000101" when "0100111011",
"10000101" when "0100111100",
"10000101" when "0100111101",
"10000101" when "0100111110",
"10000101" when "0100111111",
"10000110" when "0101000000",
"10000110" when "0101000001",
"10000110" when "0101000010",
"10000110" when "0101000011",
"10000110" when "0101000100",
"10000110" when "0101000101",
"10000110" when "0101000110",
"10000110" when "0101000111",
"10000110" when "0101001000",
"10000110" when "0101001001",
"10000110" when "0101001010",
"10000110" when "0101001011",
"10000110" when "0101001100",
"10000110" when "0101001101",
"10000110" when "0101001110",
"10000110" when "0101001111",
"10000110" when "0101010000",
"10000110" when "0101010001",
"10000110" when "0101010010",
"10000110" when "0101010011",
"10000110" when "0101010100",
"10000110" when "0101010101",
"10000110" when "0101010110",
"10000110" when "0101010111",
"10000110" when "0101011000",
"10000110" when "0101011001",
"10000110" when "0101011010",
"10000110" when "0101011011",
"10000110" when "0101011100",
"10000110" when "0101011101",
"10000110" when "0101011110",
"10000110" when "0101011111",
"10000110" when "0101100000",
"10000110" when "0101100001",
"10000110" when "0101100010",
"10000110" when "0101100011",
"10000110" when "0101100100",
"10000110" when "0101100101",
"10000110" when "0101100110",
"10000110" when "0101100111",
"10000110" when "0101101000",
"10000110" when "0101101001",
"10000110" when "0101101010",
"10000110" when "0101101011",
"10000110" when "0101101100",
"10000110" when "0101101101",
"10000110" when "0101101110",
"10000110" when "0101101111",
"10000110" when "0101110000",
"10000110" when "0101110001",
"10000110" when "0101110010",
"10000110" when "0101110011",
"10000110" when "0101110100",
"10000110" when "0101110101",
"10000110" when "0101110110",
"10000110" when "0101110111",
"10000110" when "0101111000",
"10000110" when "0101111001",
"10000110" when "0101111010",
"10000110" when "0101111011",
"10000110" when "0101111100",
"10000110" when "0101111101",
"10000110" when "0101111110",
"10000110" when "0101111111",
"10000111" when "0110000000",
"10000111" when "0110000001",
"10000111" when "0110000010",
"10000111" when "0110000011",
"10000111" when "0110000100",
"10000111" when "0110000101",
"10000111" when "0110000110",
"10000111" when "0110000111",
"10000111" when "0110001000",
"10000111" when "0110001001",
"10000111" when "0110001010",
"10000111" when "0110001011",
"10000111" when "0110001100",
"10000111" when "0110001101",
"10000111" when "0110001110",
"10000111" when "0110001111",
"10000111" when "0110010000",
"10000111" when "0110010001",
"10000111" when "0110010010",
"10000111" when "0110010011",
"10000111" when "0110010100",
"10000111" when "0110010101",
"10000111" when "0110010110",
"10000111" when "0110010111",
"10000111" when "0110011000",
"10000111" when "0110011001",
"10000111" when "0110011010",
"10000111" when "0110011011",
"10000111" when "0110011100",
"10000111" when "0110011101",
"10000111" when "0110011110",
"10000111" when "0110011111",
"10000111" when "0110100000",
"10000111" when "0110100001",
"10000111" when "0110100010",
"10000111" when "0110100011",
"10000111" when "0110100100",
"10000111" when "0110100101",
"10000111" when "0110100110",
"10000111" when "0110100111",
"10000111" when "0110101000",
"10000111" when "0110101001",
"10000111" when "0110101010",
"10000111" when "0110101011",
"10000111" when "0110101100",
"10000111" when "0110101101",
"10000111" when "0110101110",
"10000111" when "0110101111",
"10000111" when "0110110000",
"10000111" when "0110110001",
"10000111" when "0110110010",
"10000111" when "0110110011",
"10000111" when "0110110100",
"10000111" when "0110110101",
"10000111" when "0110110110",
"10000111" when "0110110111",
"10000111" when "0110111000",
"10000111" when "0110111001",
"10000111" when "0110111010",
"10000111" when "0110111011",
"10000111" when "0110111100",
"10000111" when "0110111101",
"10000111" when "0110111110",
"10000111" when "0110111111",
"10000111" when "0111000000",
"10000111" when "0111000001",
"10000111" when "0111000010",
"10000111" when "0111000011",
"10000111" when "0111000100",
"10000111" when "0111000101",
"10000111" when "0111000110",
"10000111" when "0111000111",
"10000111" when "0111001000",
"10000111" when "0111001001",
"10000111" when "0111001010",
"10000111" when "0111001011",
"10000111" when "0111001100",
"10000111" when "0111001101",
"10000111" when "0111001110",
"10000111" when "0111001111",
"10000111" when "0111010000",
"10000111" when "0111010001",
"10000111" when "0111010010",
"10000111" when "0111010011",
"10000111" when "0111010100",
"10000111" when "0111010101",
"10000111" when "0111010110",
"10000111" when "0111010111",
"10000111" when "0111011000",
"10000111" when "0111011001",
"10000111" when "0111011010",
"10000111" when "0111011011",
"10000111" when "0111011100",
"10000111" when "0111011101",
"10000111" when "0111011110",
"10000111" when "0111011111",
"10000111" when "0111100000",
"10000111" when "0111100001",
"10000111" when "0111100010",
"10000111" when "0111100011",
"10000111" when "0111100100",
"10000111" when "0111100101",
"10000111" when "0111100110",
"10000111" when "0111100111",
"10000111" when "0111101000",
"10000111" when "0111101001",
"10000111" when "0111101010",
"10000111" when "0111101011",
"10000111" when "0111101100",
"10000111" when "0111101101",
"10000111" when "0111101110",
"10000111" when "0111101111",
"10000111" when "0111110000",
"10000111" when "0111110001",
"10000111" when "0111110010",
"10000111" when "0111110011",
"10000111" when "0111110100",
"10000111" when "0111110101",
"10000111" when "0111110110",
"10000111" when "0111110111",
"10000111" when "0111111000",
"10000111" when "0111111001",
"10000111" when "0111111010",
"10000111" when "0111111011",
"10000111" when "0111111100",
"10000111" when "0111111101",
"10000111" when "0111111110",
"10000111" when "0111111111",
"10011111" when "1000000000",
"10010000" when "1000000001",
"10010001" when "1000000010",
"10010001" when "1000000011",
"10010010" when "1000000100",
"10010010" when "1000000101",
"10010010" when "1000000110",
"10010010" when "1000000111",
"10010011" when "1000001000",
"10010011" when "1000001001",
"10010011" when "1000001010",
"10010011" when "1000001011",
"10010011" when "1000001100",
"10010011" when "1000001101",
"10010011" when "1000001110",
"10010011" when "1000001111",
"10010100" when "1000010000",
"10010100" when "1000010001",
"10010100" when "1000010010",
"10010100" when "1000010011",
"10010100" when "1000010100",
"10010100" when "1000010101",
"10010100" when "1000010110",
"10010100" when "1000010111",
"10010100" when "1000011000",
"10010100" when "1000011001",
"10010100" when "1000011010",
"10010100" when "1000011011",
"10010100" when "1000011100",
"10010100" when "1000011101",
"10010100" when "1000011110",
"10010100" when "1000011111",
"10010101" when "1000100000",
"10010101" when "1000100001",
"10010101" when "1000100010",
"10010101" when "1000100011",
"10010101" when "1000100100",
"10010101" when "1000100101",
"10010101" when "1000100110",
"10010101" when "1000100111",
"10010101" when "1000101000",
"10010101" when "1000101001",
"10010101" when "1000101010",
"10010101" when "1000101011",
"10010101" when "1000101100",
"10010101" when "1000101101",
"10010101" when "1000101110",
"10010101" when "1000101111",
"10010101" when "1000110000",
"10010101" when "1000110001",
"10010101" when "1000110010",
"10010101" when "1000110011",
"10010101" when "1000110100",
"10010101" when "1000110101",
"10010101" when "1000110110",
"10010101" when "1000110111",
"10010101" when "1000111000",
"10010101" when "1000111001",
"10010101" when "1000111010",
"10010101" when "1000111011",
"10010101" when "1000111100",
"10010101" when "1000111101",
"10010101" when "1000111110",
"10010101" when "1000111111",
"10010110" when "1001000000",
"10010110" when "1001000001",
"10010110" when "1001000010",
"10010110" when "1001000011",
"10010110" when "1001000100",
"10010110" when "1001000101",
"10010110" when "1001000110",
"10010110" when "1001000111",
"10010110" when "1001001000",
"10010110" when "1001001001",
"10010110" when "1001001010",
"10010110" when "1001001011",
"10010110" when "1001001100",
"10010110" when "1001001101",
"10010110" when "1001001110",
"10010110" when "1001001111",
"10010110" when "1001010000",
"10010110" when "1001010001",
"10010110" when "1001010010",
"10010110" when "1001010011",
"10010110" when "1001010100",
"10010110" when "1001010101",
"10010110" when "1001010110",
"10010110" when "1001010111",
"10010110" when "1001011000",
"10010110" when "1001011001",
"10010110" when "1001011010",
"10010110" when "1001011011",
"10010110" when "1001011100",
"10010110" when "1001011101",
"10010110" when "1001011110",
"10010110" when "1001011111",
"10010110" when "1001100000",
"10010110" when "1001100001",
"10010110" when "1001100010",
"10010110" when "1001100011",
"10010110" when "1001100100",
"10010110" when "1001100101",
"10010110" when "1001100110",
"10010110" when "1001100111",
"10010110" when "1001101000",
"10010110" when "1001101001",
"10010110" when "1001101010",
"10010110" when "1001101011",
"10010110" when "1001101100",
"10010110" when "1001101101",
"10010110" when "1001101110",
"10010110" when "1001101111",
"10010110" when "1001110000",
"10010110" when "1001110001",
"10010110" when "1001110010",
"10010110" when "1001110011",
"10010110" when "1001110100",
"10010110" when "1001110101",
"10010110" when "1001110110",
"10010110" when "1001110111",
"10010110" when "1001111000",
"10010110" when "1001111001",
"10010110" when "1001111010",
"10010110" when "1001111011",
"10010110" when "1001111100",
"10010110" when "1001111101",
"10010110" when "1001111110",
"10010110" when "1001111111",
"10010111" when "1010000000",
"10010111" when "1010000001",
"10010111" when "1010000010",
"10010111" when "1010000011",
"10010111" when "1010000100",
"10010111" when "1010000101",
"10010111" when "1010000110",
"10010111" when "1010000111",
"10010111" when "1010001000",
"10010111" when "1010001001",
"10010111" when "1010001010",
"10010111" when "1010001011",
"10010111" when "1010001100",
"10010111" when "1010001101",
"10010111" when "1010001110",
"10010111" when "1010001111",
"10010111" when "1010010000",
"10010111" when "1010010001",
"10010111" when "1010010010",
"10010111" when "1010010011",
"10010111" when "1010010100",
"10010111" when "1010010101",
"10010111" when "1010010110",
"10010111" when "1010010111",
"10010111" when "1010011000",
"10010111" when "1010011001",
"10010111" when "1010011010",
"10010111" when "1010011011",
"10010111" when "1010011100",
"10010111" when "1010011101",
"10010111" when "1010011110",
"10010111" when "1010011111",
"10010111" when "1010100000",
"10010111" when "1010100001",
"10010111" when "1010100010",
"10010111" when "1010100011",
"10010111" when "1010100100",
"10010111" when "1010100101",
"10010111" when "1010100110",
"10010111" when "1010100111",
"10010111" when "1010101000",
"10010111" when "1010101001",
"10010111" when "1010101010",
"10010111" when "1010101011",
"10010111" when "1010101100",
"10010111" when "1010101101",
"10010111" when "1010101110",
"10010111" when "1010101111",
"10010111" when "1010110000",
"10010111" when "1010110001",
"10010111" when "1010110010",
"10010111" when "1010110011",
"10010111" when "1010110100",
"10010111" when "1010110101",
"10010111" when "1010110110",
"10010111" when "1010110111",
"10010111" when "1010111000",
"10010111" when "1010111001",
"10010111" when "1010111010",
"10010111" when "1010111011",
"10010111" when "1010111100",
"10010111" when "1010111101",
"10010111" when "1010111110",
"10010111" when "1010111111",
"10010111" when "1011000000",
"10010111" when "1011000001",
"10010111" when "1011000010",
"10010111" when "1011000011",
"10010111" when "1011000100",
"10010111" when "1011000101",
"10010111" when "1011000110",
"10010111" when "1011000111",
"10010111" when "1011001000",
"10010111" when "1011001001",
"10010111" when "1011001010",
"10010111" when "1011001011",
"10010111" when "1011001100",
"10010111" when "1011001101",
"10010111" when "1011001110",
"10010111" when "1011001111",
"10010111" when "1011010000",
"10010111" when "1011010001",
"10010111" when "1011010010",
"10010111" when "1011010011",
"10010111" when "1011010100",
"10010111" when "1011010101",
"10010111" when "1011010110",
"10010111" when "1011010111",
"10010111" when "1011011000",
"10010111" when "1011011001",
"10010111" when "1011011010",
"10010111" when "1011011011",
"10010111" when "1011011100",
"10010111" when "1011011101",
"10010111" when "1011011110",
"10010111" when "1011011111",
"10010111" when "1011100000",
"10010111" when "1011100001",
"10010111" when "1011100010",
"10010111" when "1011100011",
"10010111" when "1011100100",
"10010111" when "1011100101",
"10010111" when "1011100110",
"10010111" when "1011100111",
"10010111" when "1011101000",
"10010111" when "1011101001",
"10010111" when "1011101010",
"10010111" when "1011101011",
"10010111" when "1011101100",
"10010111" when "1011101101",
"10010111" when "1011101110",
"10010111" when "1011101111",
"10010111" when "1011110000",
"10010111" when "1011110001",
"10010111" when "1011110010",
"10010111" when "1011110011",
"10010111" when "1011110100",
"10010111" when "1011110101",
"10010111" when "1011110110",
"10010111" when "1011110111",
"10010111" when "1011111000",
"10010111" when "1011111001",
"10010111" when "1011111010",
"10010111" when "1011111011",
"10010111" when "1011111100",
"10010111" when "1011111101",
"10010111" when "1011111110",
"10010111" when "1011111111",
"10011000" when "1100000000",
"10011000" when "1100000001",
"10011000" when "1100000010",
"10011000" when "1100000011",
"10011000" when "1100000100",
"10011000" when "1100000101",
"10011000" when "1100000110",
"10011000" when "1100000111",
"10011000" when "1100001000",
"10011000" when "1100001001",
"10011000" when "1100001010",
"10011000" when "1100001011",
"10011000" when "1100001100",
"10011000" when "1100001101",
"10011000" when "1100001110",
"10011000" when "1100001111",
"10011000" when "1100010000",
"10011000" when "1100010001",
"10011000" when "1100010010",
"10011000" when "1100010011",
"10011000" when "1100010100",
"10011000" when "1100010101",
"10011000" when "1100010110",
"10011000" when "1100010111",
"10011000" when "1100011000",
"10011000" when "1100011001",
"10011000" when "1100011010",
"10011000" when "1100011011",
"10011000" when "1100011100",
"10011000" when "1100011101",
"10011000" when "1100011110",
"10011000" when "1100011111",
"10011000" when "1100100000",
"10011000" when "1100100001",
"10011000" when "1100100010",
"10011000" when "1100100011",
"10011000" when "1100100100",
"10011000" when "1100100101",
"10011000" when "1100100110",
"10011000" when "1100100111",
"10011000" when "1100101000",
"10011000" when "1100101001",
"10011000" when "1100101010",
"10011000" when "1100101011",
"10011000" when "1100101100",
"10011000" when "1100101101",
"10011000" when "1100101110",
"10011000" when "1100101111",
"10011000" when "1100110000",
"10011000" when "1100110001",
"10011000" when "1100110010",
"10011000" when "1100110011",
"10011000" when "1100110100",
"10011000" when "1100110101",
"10011000" when "1100110110",
"10011000" when "1100110111",
"10011000" when "1100111000",
"10011000" when "1100111001",
"10011000" when "1100111010",
"10011000" when "1100111011",
"10011000" when "1100111100",
"10011000" when "1100111101",
"10011000" when "1100111110",
"10011000" when "1100111111",
"10011000" when "1101000000",
"10011000" when "1101000001",
"10011000" when "1101000010",
"10011000" when "1101000011",
"10011000" when "1101000100",
"10011000" when "1101000101",
"10011000" when "1101000110",
"10011000" when "1101000111",
"10011000" when "1101001000",
"10011000" when "1101001001",
"10011000" when "1101001010",
"10011000" when "1101001011",
"10011000" when "1101001100",
"10011000" when "1101001101",
"10011000" when "1101001110",
"10011000" when "1101001111",
"10011000" when "1101010000",
"10011000" when "1101010001",
"10011000" when "1101010010",
"10011000" when "1101010011",
"10011000" when "1101010100",
"10011000" when "1101010101",
"10011000" when "1101010110",
"10011000" when "1101010111",
"10011000" when "1101011000",
"10011000" when "1101011001",
"10011000" when "1101011010",
"10011000" when "1101011011",
"10011000" when "1101011100",
"10011000" when "1101011101",
"10011000" when "1101011110",
"10011000" when "1101011111",
"10011000" when "1101100000",
"10011000" when "1101100001",
"10011000" when "1101100010",
"10011000" when "1101100011",
"10011000" when "1101100100",
"10011000" when "1101100101",
"10011000" when "1101100110",
"10011000" when "1101100111",
"10011000" when "1101101000",
"10011000" when "1101101001",
"10011000" when "1101101010",
"10011000" when "1101101011",
"10011000" when "1101101100",
"10011000" when "1101101101",
"10011000" when "1101101110",
"10011000" when "1101101111",
"10011000" when "1101110000",
"10011000" when "1101110001",
"10011000" when "1101110010",
"10011000" when "1101110011",
"10011000" when "1101110100",
"10011000" when "1101110101",
"10011000" when "1101110110",
"10011000" when "1101110111",
"10011000" when "1101111000",
"10011000" when "1101111001",
"10011000" when "1101111010",
"10011000" when "1101111011",
"10011000" when "1101111100",
"10011000" when "1101111101",
"10011000" when "1101111110",
"10011000" when "1101111111",
"10011000" when "1110000000",
"10011000" when "1110000001",
"10011000" when "1110000010",
"10011000" when "1110000011",
"10011000" when "1110000100",
"10011000" when "1110000101",
"10011000" when "1110000110",
"10011000" when "1110000111",
"10011000" when "1110001000",
"10011000" when "1110001001",
"10011000" when "1110001010",
"10011000" when "1110001011",
"10011000" when "1110001100",
"10011000" when "1110001101",
"10011000" when "1110001110",
"10011000" when "1110001111",
"10011000" when "1110010000",
"10011000" when "1110010001",
"10011000" when "1110010010",
"10011000" when "1110010011",
"10011000" when "1110010100",
"10011000" when "1110010101",
"10011000" when "1110010110",
"10011000" when "1110010111",
"10011000" when "1110011000",
"10011000" when "1110011001",
"10011000" when "1110011010",
"10011000" when "1110011011",
"10011000" when "1110011100",
"10011000" when "1110011101",
"10011000" when "1110011110",
"10011000" when "1110011111",
"10011000" when "1110100000",
"10011000" when "1110100001",
"10011000" when "1110100010",
"10011000" when "1110100011",
"10011000" when "1110100100",
"10011000" when "1110100101",
"10011000" when "1110100110",
"10011000" when "1110100111",
"10011000" when "1110101000",
"10011000" when "1110101001",
"10011000" when "1110101010",
"10011000" when "1110101011",
"10011000" when "1110101100",
"10011000" when "1110101101",
"10011000" when "1110101110",
"10011000" when "1110101111",
"10011000" when "1110110000",
"10011000" when "1110110001",
"10011000" when "1110110010",
"10011000" when "1110110011",
"10011000" when "1110110100",
"10011000" when "1110110101",
"10011000" when "1110110110",
"10011000" when "1110110111",
"10011000" when "1110111000",
"10011000" when "1110111001",
"10011000" when "1110111010",
"10011000" when "1110111011",
"10011000" when "1110111100",
"10011000" when "1110111101",
"10011000" when "1110111110",
"10011000" when "1110111111",
"10011000" when "1111000000",
"10011000" when "1111000001",
"10011000" when "1111000010",
"10011000" when "1111000011",
"10011000" when "1111000100",
"10011000" when "1111000101",
"10011000" when "1111000110",
"10011000" when "1111000111",
"10011000" when "1111001000",
"10011000" when "1111001001",
"10011000" when "1111001010",
"10011000" when "1111001011",
"10011000" when "1111001100",
"10011000" when "1111001101",
"10011000" when "1111001110",
"10011000" when "1111001111",
"10011000" when "1111010000",
"10011000" when "1111010001",
"10011000" when "1111010010",
"10011000" when "1111010011",
"10011000" when "1111010100",
"10011000" when "1111010101",
"10011000" when "1111010110",
"10011000" when "1111010111",
"10011000" when "1111011000",
"10011000" when "1111011001",
"10011000" when "1111011010",
"10011000" when "1111011011",
"10011000" when "1111011100",
"10011000" when "1111011101",
"10011000" when "1111011110",
"10011000" when "1111011111",
"10011000" when "1111100000",
"10011000" when "1111100001",
"10011000" when "1111100010",
"10011000" when "1111100011",
"10011000" when "1111100100",
"10011000" when "1111100101",
"10011000" when "1111100110",
"10011000" when "1111100111",
"10011000" when "1111101000",
"10011000" when "1111101001",
"10011000" when "1111101010",
"10011000" when "1111101011",
"10011000" when "1111101100",
"10011000" when "1111101101",
"10011000" when "1111101110",
"10011000" when "1111101111",
"10011000" when "1111110000",
"10011000" when "1111110001",
"10011000" when "1111110010",
"10011000" when "1111110011",
"10011000" when "1111110100",
"10011000" when "1111110101",
"10011000" when "1111110110",
"10011000" when "1111110111",
"10011000" when "1111111000",
"10011000" when "1111111001",
"10011000" when "1111111010",
"10011000" when "1111111011",
"10011000" when "1111111100",
"10011000" when "1111111101",
"10011000" when "1111111110",
"10011000" when others;
					
	
	fst <= both(7 downto 4);
	snd <= both(3 downto 0);

END table_arch;