library verilog;
use verilog.vl_types.all;
entity eq2_vlg_vec_tst is
end eq2_vlg_vec_tst;
