library verilog;
use verilog.vl_types.all;
entity eq2_vlg_check_tst is
    port(
        aeqb            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end eq2_vlg_check_tst;
