library verilog;
use verilog.vl_types.all;
entity zero_top_vlg_vec_tst is
end zero_top_vlg_vec_tst;
